//external port declaration and create a module
module half_adder(a,b,sum,carry);

//port direction
output a,b; //input
output sum,carry;//output
//reg sum,carry;//output
  //updated logic 
endmodule
